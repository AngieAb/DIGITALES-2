library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all; 

Entity Ale_0a5 is 

Port(Clock,Reset,Enable,Load : 	IN std_logic;
	Q: Out std_logic_vector (2 downto 0));
End Ale_0a5;

Architecture sol of Ale_0a5 is 
Begin 
end sol;
