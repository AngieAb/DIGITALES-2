library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Bin_Dec_led is
port (A: in std_logic_vector (2 downto 0);
      B: out std_logic_vector (4 downto 0));
        end Bin_Dec_led;
architecture solution of Bin_Dec_led is
begin
end solution;
